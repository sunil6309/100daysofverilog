module bufi(input en,
	input a,
	output b);
assign b= en&a;
endmodule
