module encoder(en,in,out);
  input en;
  input[7:0]in;
  output reg[2:0]out;
  if(~en)
    out<=3'd0;
  else
    begin
      case(in)
        8'b0000_0001:out=3'd0;
        8'b0000_0010:out=3'd1;
        8'b0000_0100:out=3'd2;
        8'b0000_1000:out=3'd3;
        8'b0001_0000:out=3'd4;
        8'b0010_0000:out=3'd5;
        8'b0100_0000:out=3'd6;
        8'b1000_0000:out=3'd7;
      endcase
    end
endmodule
